/*  This file is part of JTFRAME.
    JTFRAME program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTFRAME program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTFRAME. If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 11-8-2022 */

module jtframe_logo #(parameter
    COLORW = 4
) (
    input        clk,
    input        pxl_cen,
    input        show_en,

    // input  [1:0] rotate, //[0] - rotate [1] - left or right

    // VGA signals coming from core
    input  [3*COLORW-1:0] rgb_in,
    input        hs,
    input        vs,
    input        lhbl,
    input        lvbl,

    // VGA signals going to video connector
    output [3*COLORW-1:0] rgb_out,

    output reg       hs_out,
    output reg       vs_out,
    output reg       lhbl_out,
    output reg       lvbl_out
);

reg  [ 8:0] hcnt=0,vcnt=0, htot=9'd256, vtot=9'd256;
reg         hsl, vsl;
wire [10:0] addr;
reg  [ 7:0] char;
reg  [ 7:0] rom[0:8*256-1];
wire        pxl;
wire [COLORW-1:0] r_in, g_in, b_in;
reg  [COLORW-1:0] r_out, g_out, b_out;

assign addr = { vcnt[7:5], hcnt[7:0] };
assign pxl  = char[ vcnt[4:2] ];
assign {r_in,g_in,b_in} = rgb_in;
assign rgb_out = { r_out, g_out, b_out };

function [COLORW-1:0] filter( input [COLORW-1:0] a );
    filter = show_en ? {COLORW{pxl}} : a;
endfunction

always @(posedge clk) if( pxl_cen ) begin
    { hs_out, vs_out }   <= { hs, vs };
    { lhbl_out, lvbl_out } <= { lhbl, lvbl };
    r_out <= filter( r_in );
    g_out <= filter( g_in );
    b_out <= filter( b_in );
end

// screen counter
always @(posedge clk) if( pxl_cen ) begin
    hsl <= hs;
    vsl <= vs;
    hcnt <= hcnt + 9'd1;
    if( hs & ~hsl ) begin
        htot <= hcnt;
        hcnt <= 0;
        if( lvbl ) vcnt <= vcnt+9'd1;
    end
    if( vs && !vsl && vcnt!=0 ) begin
        vtot <= vcnt;
    end
end

always @(posedge clk) begin
    char <= rom[addr];
end

initial begin
    rom[   0 ] = 8'h00;
    rom[   1 ] = 8'h00;
    rom[   2 ] = 8'h00;
    rom[   3 ] = 8'h00;
    rom[   4 ] = 8'h00;
    rom[   5 ] = 8'h00;
    rom[   6 ] = 8'h00;
    rom[   7 ] = 8'h00;
    rom[   8 ] = 8'h00;
    rom[   9 ] = 8'h00;
    rom[  10 ] = 8'h00;
    rom[  11 ] = 8'h00;
    rom[  12 ] = 8'h00;
    rom[  13 ] = 8'h00;
    rom[  14 ] = 8'h00;
    rom[  15 ] = 8'h00;
    rom[  16 ] = 8'h00;
    rom[  17 ] = 8'h00;
    rom[  18 ] = 8'h00;
    rom[  19 ] = 8'h00;
    rom[  20 ] = 8'h00;
    rom[  21 ] = 8'h00;
    rom[  22 ] = 8'h00;
    rom[  23 ] = 8'h00;
    rom[  24 ] = 8'h00;
    rom[  25 ] = 8'h00;
    rom[  26 ] = 8'h00;
    rom[  27 ] = 8'h00;
    rom[  28 ] = 8'h00;
    rom[  29 ] = 8'h00;
    rom[  30 ] = 8'h00;
    rom[  31 ] = 8'h00;
    rom[  32 ] = 8'h00;
    rom[  33 ] = 8'h00;
    rom[  34 ] = 8'h00;
    rom[  35 ] = 8'h00;
    rom[  36 ] = 8'h00;
    rom[  37 ] = 8'h00;
    rom[  38 ] = 8'h00;
    rom[  39 ] = 8'h00;
    rom[  40 ] = 8'h00;
    rom[  41 ] = 8'h00;
    rom[  42 ] = 8'h00;
    rom[  43 ] = 8'h00;
    rom[  44 ] = 8'h00;
    rom[  45 ] = 8'h00;
    rom[  46 ] = 8'h00;
    rom[  47 ] = 8'h00;
    rom[  48 ] = 8'h00;
    rom[  49 ] = 8'h00;
    rom[  50 ] = 8'h00;
    rom[  51 ] = 8'h00;
    rom[  52 ] = 8'h00;
    rom[  53 ] = 8'h00;
    rom[  54 ] = 8'h00;
    rom[  55 ] = 8'h00;
    rom[  56 ] = 8'h00;
    rom[  57 ] = 8'h00;
    rom[  58 ] = 8'h00;
    rom[  59 ] = 8'h00;
    rom[  60 ] = 8'h00;
    rom[  61 ] = 8'h00;
    rom[  62 ] = 8'h00;
    rom[  63 ] = 8'h00;
    rom[  64 ] = 8'h00;
    rom[  65 ] = 8'h00;
    rom[  66 ] = 8'h00;
    rom[  67 ] = 8'h00;
    rom[  68 ] = 8'h00;
    rom[  69 ] = 8'h00;
    rom[  70 ] = 8'h00;
    rom[  71 ] = 8'h00;
    rom[  72 ] = 8'h00;
    rom[  73 ] = 8'h00;
    rom[  74 ] = 8'h00;
    rom[  75 ] = 8'h00;
    rom[  76 ] = 8'h00;
    rom[  77 ] = 8'h00;
    rom[  78 ] = 8'h00;
    rom[  79 ] = 8'h00;
    rom[  80 ] = 8'h00;
    rom[  81 ] = 8'h00;
    rom[  82 ] = 8'h00;
    rom[  83 ] = 8'h00;
    rom[  84 ] = 8'h00;
    rom[  85 ] = 8'h00;
    rom[  86 ] = 8'h00;
    rom[  87 ] = 8'h00;
    rom[  88 ] = 8'h00;
    rom[  89 ] = 8'h00;
    rom[  90 ] = 8'h00;
    rom[  91 ] = 8'h00;
    rom[  92 ] = 8'h00;
    rom[  93 ] = 8'h00;
    rom[  94 ] = 8'h00;
    rom[  95 ] = 8'h00;
    rom[  96 ] = 8'h00;
    rom[  97 ] = 8'h00;
    rom[  98 ] = 8'h00;
    rom[  99 ] = 8'h00;
    rom[ 100 ] = 8'h00;
    rom[ 101 ] = 8'h00;
    rom[ 102 ] = 8'h00;
    rom[ 103 ] = 8'h00;
    rom[ 104 ] = 8'h00;
    rom[ 105 ] = 8'h00;
    rom[ 106 ] = 8'h00;
    rom[ 107 ] = 8'h00;
    rom[ 108 ] = 8'h00;
    rom[ 109 ] = 8'h00;
    rom[ 110 ] = 8'h00;
    rom[ 111 ] = 8'h00;
    rom[ 112 ] = 8'h00;
    rom[ 113 ] = 8'h00;
    rom[ 114 ] = 8'h00;
    rom[ 115 ] = 8'h00;
    rom[ 116 ] = 8'h00;
    rom[ 117 ] = 8'h00;
    rom[ 118 ] = 8'h00;
    rom[ 119 ] = 8'h00;
    rom[ 120 ] = 8'h00;
    rom[ 121 ] = 8'h00;
    rom[ 122 ] = 8'h00;
    rom[ 123 ] = 8'h00;
    rom[ 124 ] = 8'h00;
    rom[ 125 ] = 8'h00;
    rom[ 126 ] = 8'h00;
    rom[ 127 ] = 8'h00;
    rom[ 128 ] = 8'h00;
    rom[ 129 ] = 8'hC0;
    rom[ 130 ] = 8'hF0;
    rom[ 131 ] = 8'hF8;
    rom[ 132 ] = 8'hFC;
    rom[ 133 ] = 8'hFC;
    rom[ 134 ] = 8'hFC;
    rom[ 135 ] = 8'hFC;
    rom[ 136 ] = 8'hFC;
    rom[ 137 ] = 8'hFC;
    rom[ 138 ] = 8'hFC;
    rom[ 139 ] = 8'hFC;
    rom[ 140 ] = 8'hFC;
    rom[ 141 ] = 8'hFC;
    rom[ 142 ] = 8'hFC;
    rom[ 143 ] = 8'hFC;
    rom[ 144 ] = 8'hFC;
    rom[ 145 ] = 8'hFC;
    rom[ 146 ] = 8'hFC;
    rom[ 147 ] = 8'hFC;
    rom[ 148 ] = 8'hFC;
    rom[ 149 ] = 8'hFC;
    rom[ 150 ] = 8'hFC;
    rom[ 151 ] = 8'hFC;
    rom[ 152 ] = 8'hFC;
    rom[ 153 ] = 8'hFC;
    rom[ 154 ] = 8'hFC;
    rom[ 155 ] = 8'hFC;
    rom[ 156 ] = 8'hFC;
    rom[ 157 ] = 8'hFC;
    rom[ 158 ] = 8'hFC;
    rom[ 159 ] = 8'hFC;
    rom[ 160 ] = 8'hF0;
    rom[ 161 ] = 8'hF0;
    rom[ 162 ] = 8'hF0;
    rom[ 163 ] = 8'hC0;
    rom[ 164 ] = 8'hC0;
    rom[ 165 ] = 8'hC0;
    rom[ 166 ] = 8'hC0;
    rom[ 167 ] = 8'hC0;
    rom[ 168 ] = 8'h00;
    rom[ 169 ] = 8'h00;
    rom[ 170 ] = 8'h00;
    rom[ 171 ] = 8'h00;
    rom[ 172 ] = 8'h00;
    rom[ 173 ] = 8'h00;
    rom[ 174 ] = 8'h00;
    rom[ 175 ] = 8'h00;
    rom[ 176 ] = 8'h00;
    rom[ 177 ] = 8'h00;
    rom[ 178 ] = 8'h00;
    rom[ 179 ] = 8'h00;
    rom[ 180 ] = 8'h00;
    rom[ 181 ] = 8'h00;
    rom[ 182 ] = 8'h00;
    rom[ 183 ] = 8'h00;
    rom[ 184 ] = 8'h00;
    rom[ 185 ] = 8'h00;
    rom[ 186 ] = 8'h00;
    rom[ 187 ] = 8'h00;
    rom[ 188 ] = 8'h00;
    rom[ 189 ] = 8'h00;
    rom[ 190 ] = 8'h00;
    rom[ 191 ] = 8'h00;
    rom[ 192 ] = 8'h00;
    rom[ 193 ] = 8'h00;
    rom[ 194 ] = 8'h00;
    rom[ 195 ] = 8'h00;
    rom[ 196 ] = 8'h00;
    rom[ 197 ] = 8'h00;
    rom[ 198 ] = 8'h00;
    rom[ 199 ] = 8'h00;
    rom[ 200 ] = 8'h00;
    rom[ 201 ] = 8'h00;
    rom[ 202 ] = 8'h00;
    rom[ 203 ] = 8'h00;
    rom[ 204 ] = 8'h00;
    rom[ 205 ] = 8'h00;
    rom[ 206 ] = 8'h00;
    rom[ 207 ] = 8'h00;
    rom[ 208 ] = 8'h00;
    rom[ 209 ] = 8'h00;
    rom[ 210 ] = 8'h00;
    rom[ 211 ] = 8'h00;
    rom[ 212 ] = 8'h00;
    rom[ 213 ] = 8'h00;
    rom[ 214 ] = 8'h00;
    rom[ 215 ] = 8'h00;
    rom[ 216 ] = 8'h00;
    rom[ 217 ] = 8'h00;
    rom[ 218 ] = 8'h00;
    rom[ 219 ] = 8'h00;
    rom[ 220 ] = 8'h00;
    rom[ 221 ] = 8'h00;
    rom[ 222 ] = 8'h00;
    rom[ 223 ] = 8'h00;
    rom[ 224 ] = 8'h00;
    rom[ 225 ] = 8'h00;
    rom[ 226 ] = 8'h00;
    rom[ 227 ] = 8'h00;
    rom[ 228 ] = 8'h00;
    rom[ 229 ] = 8'h00;
    rom[ 230 ] = 8'h00;
    rom[ 231 ] = 8'h00;
    rom[ 232 ] = 8'h00;
    rom[ 233 ] = 8'h00;
    rom[ 234 ] = 8'h00;
    rom[ 235 ] = 8'h00;
    rom[ 236 ] = 8'h00;
    rom[ 237 ] = 8'h00;
    rom[ 238 ] = 8'h00;
    rom[ 239 ] = 8'h00;
    rom[ 240 ] = 8'h00;
    rom[ 241 ] = 8'h00;
    rom[ 242 ] = 8'h00;
    rom[ 243 ] = 8'h00;
    rom[ 244 ] = 8'h00;
    rom[ 245 ] = 8'h00;
    rom[ 246 ] = 8'h00;
    rom[ 247 ] = 8'h00;
    rom[ 248 ] = 8'h00;
    rom[ 249 ] = 8'h00;
    rom[ 250 ] = 8'h00;
    rom[ 251 ] = 8'h00;
    rom[ 252 ] = 8'h00;
    rom[ 253 ] = 8'h00;
    rom[ 254 ] = 8'h00;
    rom[ 255 ] = 8'h00;
    rom[ 256 ] = 8'h00;
    rom[ 257 ] = 8'h00;
    rom[ 258 ] = 8'h00;
    rom[ 259 ] = 8'h00;
    rom[ 260 ] = 8'h00;
    rom[ 261 ] = 8'h00;
    rom[ 262 ] = 8'h00;
    rom[ 263 ] = 8'h00;
    rom[ 264 ] = 8'h00;
    rom[ 265 ] = 8'h00;
    rom[ 266 ] = 8'h00;
    rom[ 267 ] = 8'h00;
    rom[ 268 ] = 8'h00;
    rom[ 269 ] = 8'h00;
    rom[ 270 ] = 8'h00;
    rom[ 271 ] = 8'h00;
    rom[ 272 ] = 8'h00;
    rom[ 273 ] = 8'h00;
    rom[ 274 ] = 8'h00;
    rom[ 275 ] = 8'h00;
    rom[ 276 ] = 8'h00;
    rom[ 277 ] = 8'h00;
    rom[ 278 ] = 8'h00;
    rom[ 279 ] = 8'h00;
    rom[ 280 ] = 8'h00;
    rom[ 281 ] = 8'h00;
    rom[ 282 ] = 8'h00;
    rom[ 283 ] = 8'h00;
    rom[ 284 ] = 8'h00;
    rom[ 285 ] = 8'h00;
    rom[ 286 ] = 8'h00;
    rom[ 287 ] = 8'h00;
    rom[ 288 ] = 8'h00;
    rom[ 289 ] = 8'h00;
    rom[ 290 ] = 8'h00;
    rom[ 291 ] = 8'h00;
    rom[ 292 ] = 8'h00;
    rom[ 293 ] = 8'h00;
    rom[ 294 ] = 8'h00;
    rom[ 295 ] = 8'h00;
    rom[ 296 ] = 8'h00;
    rom[ 297 ] = 8'h00;
    rom[ 298 ] = 8'h00;
    rom[ 299 ] = 8'h00;
    rom[ 300 ] = 8'h00;
    rom[ 301 ] = 8'h00;
    rom[ 302 ] = 8'h00;
    rom[ 303 ] = 8'h00;
    rom[ 304 ] = 8'h00;
    rom[ 305 ] = 8'h00;
    rom[ 306 ] = 8'h00;
    rom[ 307 ] = 8'h00;
    rom[ 308 ] = 8'h00;
    rom[ 309 ] = 8'h00;
    rom[ 310 ] = 8'h00;
    rom[ 311 ] = 8'h00;
    rom[ 312 ] = 8'h00;
    rom[ 313 ] = 8'h00;
    rom[ 314 ] = 8'h00;
    rom[ 315 ] = 8'h00;
    rom[ 316 ] = 8'h00;
    rom[ 317 ] = 8'h00;
    rom[ 318 ] = 8'h00;
    rom[ 319 ] = 8'h00;
    rom[ 320 ] = 8'h00;
    rom[ 321 ] = 8'h00;
    rom[ 322 ] = 8'h00;
    rom[ 323 ] = 8'h00;
    rom[ 324 ] = 8'h00;
    rom[ 325 ] = 8'h00;
    rom[ 326 ] = 8'h00;
    rom[ 327 ] = 8'h00;
    rom[ 328 ] = 8'h00;
    rom[ 329 ] = 8'h00;
    rom[ 330 ] = 8'h00;
    rom[ 331 ] = 8'h00;
    rom[ 332 ] = 8'h00;
    rom[ 333 ] = 8'h00;
    rom[ 334 ] = 8'h00;
    rom[ 335 ] = 8'h00;
    rom[ 336 ] = 8'h00;
    rom[ 337 ] = 8'h00;
    rom[ 338 ] = 8'h00;
    rom[ 339 ] = 8'h00;
    rom[ 340 ] = 8'h00;
    rom[ 341 ] = 8'h00;
    rom[ 342 ] = 8'h00;
    rom[ 343 ] = 8'h00;
    rom[ 344 ] = 8'h00;
    rom[ 345 ] = 8'h00;
    rom[ 346 ] = 8'h00;
    rom[ 347 ] = 8'h00;
    rom[ 348 ] = 8'h00;
    rom[ 349 ] = 8'h00;
    rom[ 350 ] = 8'h00;
    rom[ 351 ] = 8'h00;
    rom[ 352 ] = 8'h00;
    rom[ 353 ] = 8'h00;
    rom[ 354 ] = 8'h00;
    rom[ 355 ] = 8'h00;
    rom[ 356 ] = 8'h00;
    rom[ 357 ] = 8'h00;
    rom[ 358 ] = 8'h00;
    rom[ 359 ] = 8'h00;
    rom[ 360 ] = 8'h00;
    rom[ 361 ] = 8'h00;
    rom[ 362 ] = 8'h80;
    rom[ 363 ] = 8'hC0;
    rom[ 364 ] = 8'hF0;
    rom[ 365 ] = 8'hF8;
    rom[ 366 ] = 8'hF8;
    rom[ 367 ] = 8'hF8;
    rom[ 368 ] = 8'hF8;
    rom[ 369 ] = 8'hF8;
    rom[ 370 ] = 8'hF8;
    rom[ 371 ] = 8'hF8;
    rom[ 372 ] = 8'hF8;
    rom[ 373 ] = 8'hF8;
    rom[ 374 ] = 8'hF8;
    rom[ 375 ] = 8'hF8;
    rom[ 376 ] = 8'hF8;
    rom[ 377 ] = 8'hF8;
    rom[ 378 ] = 8'hF8;
    rom[ 379 ] = 8'hF8;
    rom[ 380 ] = 8'hF8;
    rom[ 381 ] = 8'hF8;
    rom[ 382 ] = 8'hF8;
    rom[ 383 ] = 8'hFC;
    rom[ 384 ] = 8'hFF;
    rom[ 385 ] = 8'hFF;
    rom[ 386 ] = 8'hFF;
    rom[ 387 ] = 8'hFF;
    rom[ 388 ] = 8'hFF;
    rom[ 389 ] = 8'hFF;
    rom[ 390 ] = 8'hFF;
    rom[ 391 ] = 8'hFF;
    rom[ 392 ] = 8'hFF;
    rom[ 393 ] = 8'hFF;
    rom[ 394 ] = 8'hFF;
    rom[ 395 ] = 8'hFF;
    rom[ 396 ] = 8'hFF;
    rom[ 397 ] = 8'hFF;
    rom[ 398 ] = 8'hFF;
    rom[ 399 ] = 8'hFF;
    rom[ 400 ] = 8'hFF;
    rom[ 401 ] = 8'hFF;
    rom[ 402 ] = 8'hFF;
    rom[ 403 ] = 8'hFF;
    rom[ 404 ] = 8'hFF;
    rom[ 405 ] = 8'hFF;
    rom[ 406 ] = 8'hFF;
    rom[ 407 ] = 8'hFF;
    rom[ 408 ] = 8'hFF;
    rom[ 409 ] = 8'hFF;
    rom[ 410 ] = 8'hFF;
    rom[ 411 ] = 8'hFF;
    rom[ 412 ] = 8'hFF;
    rom[ 413 ] = 8'hFF;
    rom[ 414 ] = 8'hFF;
    rom[ 415 ] = 8'hFF;
    rom[ 416 ] = 8'hFF;
    rom[ 417 ] = 8'hFF;
    rom[ 418 ] = 8'hFF;
    rom[ 419 ] = 8'hFF;
    rom[ 420 ] = 8'hFF;
    rom[ 421 ] = 8'hFF;
    rom[ 422 ] = 8'hF9;
    rom[ 423 ] = 8'hF8;
    rom[ 424 ] = 8'hF8;
    rom[ 425 ] = 8'hF8;
    rom[ 426 ] = 8'hF8;
    rom[ 427 ] = 8'hF8;
    rom[ 428 ] = 8'hF8;
    rom[ 429 ] = 8'hF8;
    rom[ 430 ] = 8'hF8;
    rom[ 431 ] = 8'hF8;
    rom[ 432 ] = 8'hF8;
    rom[ 433 ] = 8'hF8;
    rom[ 434 ] = 8'hF8;
    rom[ 435 ] = 8'hF8;
    rom[ 436 ] = 8'hF8;
    rom[ 437 ] = 8'hF8;
    rom[ 438 ] = 8'hF8;
    rom[ 439 ] = 8'hF8;
    rom[ 440 ] = 8'hF8;
    rom[ 441 ] = 8'hF8;
    rom[ 442 ] = 8'hF8;
    rom[ 443 ] = 8'hF8;
    rom[ 444 ] = 8'hF8;
    rom[ 445 ] = 8'hF8;
    rom[ 446 ] = 8'hF8;
    rom[ 447 ] = 8'hF8;
    rom[ 448 ] = 8'hF8;
    rom[ 449 ] = 8'hF8;
    rom[ 450 ] = 8'hF8;
    rom[ 451 ] = 8'hF8;
    rom[ 452 ] = 8'hF8;
    rom[ 453 ] = 8'hF8;
    rom[ 454 ] = 8'hF8;
    rom[ 455 ] = 8'hF8;
    rom[ 456 ] = 8'hF8;
    rom[ 457 ] = 8'hF8;
    rom[ 458 ] = 8'hF8;
    rom[ 459 ] = 8'hF8;
    rom[ 460 ] = 8'hF8;
    rom[ 461 ] = 8'hF8;
    rom[ 462 ] = 8'hF8;
    rom[ 463 ] = 8'hF8;
    rom[ 464 ] = 8'hF8;
    rom[ 465 ] = 8'hF8;
    rom[ 466 ] = 8'hF8;
    rom[ 467 ] = 8'hF8;
    rom[ 468 ] = 8'hF8;
    rom[ 469 ] = 8'hF8;
    rom[ 470 ] = 8'hF8;
    rom[ 471 ] = 8'hF8;
    rom[ 472 ] = 8'hF8;
    rom[ 473 ] = 8'hF8;
    rom[ 474 ] = 8'hF8;
    rom[ 475 ] = 8'hF8;
    rom[ 476 ] = 8'hF8;
    rom[ 477 ] = 8'hF8;
    rom[ 478 ] = 8'hF8;
    rom[ 479 ] = 8'hF8;
    rom[ 480 ] = 8'hF8;
    rom[ 481 ] = 8'hF8;
    rom[ 482 ] = 8'hF8;
    rom[ 483 ] = 8'hF8;
    rom[ 484 ] = 8'hF8;
    rom[ 485 ] = 8'hF8;
    rom[ 486 ] = 8'hF8;
    rom[ 487 ] = 8'hF8;
    rom[ 488 ] = 8'hF8;
    rom[ 489 ] = 8'hF8;
    rom[ 490 ] = 8'hF8;
    rom[ 491 ] = 8'hF8;
    rom[ 492 ] = 8'hF8;
    rom[ 493 ] = 8'hF8;
    rom[ 494 ] = 8'hF8;
    rom[ 495 ] = 8'hF8;
    rom[ 496 ] = 8'hF8;
    rom[ 497 ] = 8'hF8;
    rom[ 498 ] = 8'hF8;
    rom[ 499 ] = 8'hF8;
    rom[ 500 ] = 8'hF8;
    rom[ 501 ] = 8'hC8;
    rom[ 502 ] = 8'hC0;
    rom[ 503 ] = 8'hC0;
    rom[ 504 ] = 8'h80;
    rom[ 505 ] = 8'h80;
    rom[ 506 ] = 8'h80;
    rom[ 507 ] = 8'h80;
    rom[ 508 ] = 8'h80;
    rom[ 509 ] = 8'h00;
    rom[ 510 ] = 8'h00;
    rom[ 511 ] = 8'h00;
    rom[ 512 ] = 8'h00;
    rom[ 513 ] = 8'h00;
    rom[ 514 ] = 8'h00;
    rom[ 515 ] = 8'h00;
    rom[ 516 ] = 8'h00;
    rom[ 517 ] = 8'h00;
    rom[ 518 ] = 8'h00;
    rom[ 519 ] = 8'h00;
    rom[ 520 ] = 8'h00;
    rom[ 521 ] = 8'h00;
    rom[ 522 ] = 8'h00;
    rom[ 523 ] = 8'h00;
    rom[ 524 ] = 8'h00;
    rom[ 525 ] = 8'h00;
    rom[ 526 ] = 8'h00;
    rom[ 527 ] = 8'h00;
    rom[ 528 ] = 8'h00;
    rom[ 529 ] = 8'h00;
    rom[ 530 ] = 8'h00;
    rom[ 531 ] = 8'h00;
    rom[ 532 ] = 8'h00;
    rom[ 533 ] = 8'h00;
    rom[ 534 ] = 8'h00;
    rom[ 535 ] = 8'h00;
    rom[ 536 ] = 8'h00;
    rom[ 537 ] = 8'h00;
    rom[ 538 ] = 8'h00;
    rom[ 539 ] = 8'h00;
    rom[ 540 ] = 8'h00;
    rom[ 541 ] = 8'h00;
    rom[ 542 ] = 8'h00;
    rom[ 543 ] = 8'h00;
    rom[ 544 ] = 8'h00;
    rom[ 545 ] = 8'h00;
    rom[ 546 ] = 8'h00;
    rom[ 547 ] = 8'h00;
    rom[ 548 ] = 8'h00;
    rom[ 549 ] = 8'h00;
    rom[ 550 ] = 8'h00;
    rom[ 551 ] = 8'h00;
    rom[ 552 ] = 8'h00;
    rom[ 553 ] = 8'h00;
    rom[ 554 ] = 8'h00;
    rom[ 555 ] = 8'h00;
    rom[ 556 ] = 8'h00;
    rom[ 557 ] = 8'h00;
    rom[ 558 ] = 8'h00;
    rom[ 559 ] = 8'h00;
    rom[ 560 ] = 8'h00;
    rom[ 561 ] = 8'h00;
    rom[ 562 ] = 8'h00;
    rom[ 563 ] = 8'h00;
    rom[ 564 ] = 8'h00;
    rom[ 565 ] = 8'h00;
    rom[ 566 ] = 8'h00;
    rom[ 567 ] = 8'h00;
    rom[ 568 ] = 8'h00;
    rom[ 569 ] = 8'h00;
    rom[ 570 ] = 8'h00;
    rom[ 571 ] = 8'h00;
    rom[ 572 ] = 8'h00;
    rom[ 573 ] = 8'h00;
    rom[ 574 ] = 8'h00;
    rom[ 575 ] = 8'h00;
    rom[ 576 ] = 8'h00;
    rom[ 577 ] = 8'h00;
    rom[ 578 ] = 8'h00;
    rom[ 579 ] = 8'h00;
    rom[ 580 ] = 8'h00;
    rom[ 581 ] = 8'h00;
    rom[ 582 ] = 8'h00;
    rom[ 583 ] = 8'h00;
    rom[ 584 ] = 8'h00;
    rom[ 585 ] = 8'h00;
    rom[ 586 ] = 8'h00;
    rom[ 587 ] = 8'h00;
    rom[ 588 ] = 8'h00;
    rom[ 589 ] = 8'h00;
    rom[ 590 ] = 8'h00;
    rom[ 591 ] = 8'h00;
    rom[ 592 ] = 8'h00;
    rom[ 593 ] = 8'h00;
    rom[ 594 ] = 8'h00;
    rom[ 595 ] = 8'h00;
    rom[ 596 ] = 8'h00;
    rom[ 597 ] = 8'h00;
    rom[ 598 ] = 8'h00;
    rom[ 599 ] = 8'h00;
    rom[ 600 ] = 8'h00;
    rom[ 601 ] = 8'h00;
    rom[ 602 ] = 8'h00;
    rom[ 603 ] = 8'h00;
    rom[ 604 ] = 8'h00;
    rom[ 605 ] = 8'h00;
    rom[ 606 ] = 8'h00;
    rom[ 607 ] = 8'h00;
    rom[ 608 ] = 8'h00;
    rom[ 609 ] = 8'h00;
    rom[ 610 ] = 8'h00;
    rom[ 611 ] = 8'h00;
    rom[ 612 ] = 8'h00;
    rom[ 613 ] = 8'h00;
    rom[ 614 ] = 8'h80;
    rom[ 615 ] = 8'hE0;
    rom[ 616 ] = 8'hF8;
    rom[ 617 ] = 8'hFE;
    rom[ 618 ] = 8'hFF;
    rom[ 619 ] = 8'hFF;
    rom[ 620 ] = 8'hFF;
    rom[ 621 ] = 8'hFF;
    rom[ 622 ] = 8'hFF;
    rom[ 623 ] = 8'hFF;
    rom[ 624 ] = 8'hFF;
    rom[ 625 ] = 8'hFF;
    rom[ 626 ] = 8'hFF;
    rom[ 627 ] = 8'hFF;
    rom[ 628 ] = 8'hFF;
    rom[ 629 ] = 8'hFF;
    rom[ 630 ] = 8'hFF;
    rom[ 631 ] = 8'hFF;
    rom[ 632 ] = 8'hFF;
    rom[ 633 ] = 8'hFF;
    rom[ 634 ] = 8'hFF;
    rom[ 635 ] = 8'hFF;
    rom[ 636 ] = 8'hFF;
    rom[ 637 ] = 8'hFF;
    rom[ 638 ] = 8'hFF;
    rom[ 639 ] = 8'hFF;
    rom[ 640 ] = 8'hFF;
    rom[ 641 ] = 8'hFF;
    rom[ 642 ] = 8'hFF;
    rom[ 643 ] = 8'hFF;
    rom[ 644 ] = 8'hFF;
    rom[ 645 ] = 8'hFF;
    rom[ 646 ] = 8'hFF;
    rom[ 647 ] = 8'hFF;
    rom[ 648 ] = 8'hFF;
    rom[ 649 ] = 8'hFF;
    rom[ 650 ] = 8'hFF;
    rom[ 651 ] = 8'hFF;
    rom[ 652 ] = 8'hFF;
    rom[ 653 ] = 8'hFF;
    rom[ 654 ] = 8'hFF;
    rom[ 655 ] = 8'hFF;
    rom[ 656 ] = 8'hFF;
    rom[ 657 ] = 8'hFF;
    rom[ 658 ] = 8'hFF;
    rom[ 659 ] = 8'hFF;
    rom[ 660 ] = 8'hFF;
    rom[ 661 ] = 8'hFF;
    rom[ 662 ] = 8'hFF;
    rom[ 663 ] = 8'hFF;
    rom[ 664 ] = 8'hFF;
    rom[ 665 ] = 8'hFF;
    rom[ 666 ] = 8'hFF;
    rom[ 667 ] = 8'hFF;
    rom[ 668 ] = 8'hFF;
    rom[ 669 ] = 8'hFF;
    rom[ 670 ] = 8'hFF;
    rom[ 671 ] = 8'hFF;
    rom[ 672 ] = 8'hFF;
    rom[ 673 ] = 8'hFF;
    rom[ 674 ] = 8'hFF;
    rom[ 675 ] = 8'hFF;
    rom[ 676 ] = 8'hFF;
    rom[ 677 ] = 8'hFF;
    rom[ 678 ] = 8'hFF;
    rom[ 679 ] = 8'hFF;
    rom[ 680 ] = 8'hFF;
    rom[ 681 ] = 8'hFF;
    rom[ 682 ] = 8'hFF;
    rom[ 683 ] = 8'hFF;
    rom[ 684 ] = 8'hFF;
    rom[ 685 ] = 8'hFF;
    rom[ 686 ] = 8'hFF;
    rom[ 687 ] = 8'hFF;
    rom[ 688 ] = 8'hFF;
    rom[ 689 ] = 8'hFF;
    rom[ 690 ] = 8'hFF;
    rom[ 691 ] = 8'hFF;
    rom[ 692 ] = 8'hFF;
    rom[ 693 ] = 8'hFF;
    rom[ 694 ] = 8'hFF;
    rom[ 695 ] = 8'hFF;
    rom[ 696 ] = 8'hFF;
    rom[ 697 ] = 8'hFF;
    rom[ 698 ] = 8'hFF;
    rom[ 699 ] = 8'hFF;
    rom[ 700 ] = 8'hFF;
    rom[ 701 ] = 8'hFF;
    rom[ 702 ] = 8'hFF;
    rom[ 703 ] = 8'hFF;
    rom[ 704 ] = 8'hFF;
    rom[ 705 ] = 8'hFF;
    rom[ 706 ] = 8'hFF;
    rom[ 707 ] = 8'hFF;
    rom[ 708 ] = 8'hFF;
    rom[ 709 ] = 8'hFF;
    rom[ 710 ] = 8'hFF;
    rom[ 711 ] = 8'hFF;
    rom[ 712 ] = 8'hFF;
    rom[ 713 ] = 8'hFF;
    rom[ 714 ] = 8'hFF;
    rom[ 715 ] = 8'hFF;
    rom[ 716 ] = 8'hFF;
    rom[ 717 ] = 8'hFF;
    rom[ 718 ] = 8'hFF;
    rom[ 719 ] = 8'hFF;
    rom[ 720 ] = 8'hFF;
    rom[ 721 ] = 8'hFF;
    rom[ 722 ] = 8'hFF;
    rom[ 723 ] = 8'hFF;
    rom[ 724 ] = 8'hFF;
    rom[ 725 ] = 8'hFF;
    rom[ 726 ] = 8'hFF;
    rom[ 727 ] = 8'hFF;
    rom[ 728 ] = 8'hFF;
    rom[ 729 ] = 8'hFF;
    rom[ 730 ] = 8'hFF;
    rom[ 731 ] = 8'hFF;
    rom[ 732 ] = 8'hFF;
    rom[ 733 ] = 8'hFF;
    rom[ 734 ] = 8'hFF;
    rom[ 735 ] = 8'hFF;
    rom[ 736 ] = 8'hFF;
    rom[ 737 ] = 8'hFF;
    rom[ 738 ] = 8'hFF;
    rom[ 739 ] = 8'hFF;
    rom[ 740 ] = 8'hFF;
    rom[ 741 ] = 8'hFF;
    rom[ 742 ] = 8'hFF;
    rom[ 743 ] = 8'hFF;
    rom[ 744 ] = 8'hFF;
    rom[ 745 ] = 8'hFF;
    rom[ 746 ] = 8'hFF;
    rom[ 747 ] = 8'hFF;
    rom[ 748 ] = 8'hFF;
    rom[ 749 ] = 8'hFF;
    rom[ 750 ] = 8'hFF;
    rom[ 751 ] = 8'hFF;
    rom[ 752 ] = 8'hFF;
    rom[ 753 ] = 8'hFF;
    rom[ 754 ] = 8'hFF;
    rom[ 755 ] = 8'hFF;
    rom[ 756 ] = 8'hFF;
    rom[ 757 ] = 8'hFF;
    rom[ 758 ] = 8'hFF;
    rom[ 759 ] = 8'hFF;
    rom[ 760 ] = 8'hFF;
    rom[ 761 ] = 8'h3F;
    rom[ 762 ] = 8'h0F;
    rom[ 763 ] = 8'h07;
    rom[ 764 ] = 8'h01;
    rom[ 765 ] = 8'h00;
    rom[ 766 ] = 8'h00;
    rom[ 767 ] = 8'h00;
    rom[ 768 ] = 8'h00;
    rom[ 769 ] = 8'h00;
    rom[ 770 ] = 8'h00;
    rom[ 771 ] = 8'h00;
    rom[ 772 ] = 8'h00;
    rom[ 773 ] = 8'h00;
    rom[ 774 ] = 8'h00;
    rom[ 775 ] = 8'h00;
    rom[ 776 ] = 8'h00;
    rom[ 777 ] = 8'h00;
    rom[ 778 ] = 8'h00;
    rom[ 779 ] = 8'h00;
    rom[ 780 ] = 8'h00;
    rom[ 781 ] = 8'h00;
    rom[ 782 ] = 8'h00;
    rom[ 783 ] = 8'h00;
    rom[ 784 ] = 8'h00;
    rom[ 785 ] = 8'h00;
    rom[ 786 ] = 8'h00;
    rom[ 787 ] = 8'h00;
    rom[ 788 ] = 8'h00;
    rom[ 789 ] = 8'h00;
    rom[ 790 ] = 8'h00;
    rom[ 791 ] = 8'h00;
    rom[ 792 ] = 8'h00;
    rom[ 793 ] = 8'h00;
    rom[ 794 ] = 8'h00;
    rom[ 795 ] = 8'h00;
    rom[ 796 ] = 8'h00;
    rom[ 797 ] = 8'h00;
    rom[ 798 ] = 8'h00;
    rom[ 799 ] = 8'h00;
    rom[ 800 ] = 8'h00;
    rom[ 801 ] = 8'h00;
    rom[ 802 ] = 8'h00;
    rom[ 803 ] = 8'h00;
    rom[ 804 ] = 8'h00;
    rom[ 805 ] = 8'h00;
    rom[ 806 ] = 8'h00;
    rom[ 807 ] = 8'h00;
    rom[ 808 ] = 8'h00;
    rom[ 809 ] = 8'h00;
    rom[ 810 ] = 8'h00;
    rom[ 811 ] = 8'h00;
    rom[ 812 ] = 8'h00;
    rom[ 813 ] = 8'h00;
    rom[ 814 ] = 8'h00;
    rom[ 815 ] = 8'h00;
    rom[ 816 ] = 8'h00;
    rom[ 817 ] = 8'h00;
    rom[ 818 ] = 8'h00;
    rom[ 819 ] = 8'h00;
    rom[ 820 ] = 8'h00;
    rom[ 821 ] = 8'h00;
    rom[ 822 ] = 8'h00;
    rom[ 823 ] = 8'h00;
    rom[ 824 ] = 8'h00;
    rom[ 825 ] = 8'h00;
    rom[ 826 ] = 8'h00;
    rom[ 827 ] = 8'h00;
    rom[ 828 ] = 8'h00;
    rom[ 829 ] = 8'h00;
    rom[ 830 ] = 8'h00;
    rom[ 831 ] = 8'h00;
    rom[ 832 ] = 8'h00;
    rom[ 833 ] = 8'h00;
    rom[ 834 ] = 8'h00;
    rom[ 835 ] = 8'h00;
    rom[ 836 ] = 8'h00;
    rom[ 837 ] = 8'h00;
    rom[ 838 ] = 8'h00;
    rom[ 839 ] = 8'h00;
    rom[ 840 ] = 8'h00;
    rom[ 841 ] = 8'h00;
    rom[ 842 ] = 8'h00;
    rom[ 843 ] = 8'h00;
    rom[ 844 ] = 8'h00;
    rom[ 845 ] = 8'h00;
    rom[ 846 ] = 8'h00;
    rom[ 847 ] = 8'h00;
    rom[ 848 ] = 8'h00;
    rom[ 849 ] = 8'h00;
    rom[ 850 ] = 8'h00;
    rom[ 851 ] = 8'h00;
    rom[ 852 ] = 8'h00;
    rom[ 853 ] = 8'h00;
    rom[ 854 ] = 8'h00;
    rom[ 855 ] = 8'h00;
    rom[ 856 ] = 8'h00;
    rom[ 857 ] = 8'h00;
    rom[ 858 ] = 8'h00;
    rom[ 859 ] = 8'h00;
    rom[ 860 ] = 8'h00;
    rom[ 861 ] = 8'h00;
    rom[ 862 ] = 8'h00;
    rom[ 863 ] = 8'h00;
    rom[ 864 ] = 8'h00;
    rom[ 865 ] = 8'h00;
    rom[ 866 ] = 8'h00;
    rom[ 867 ] = 8'h00;
    rom[ 868 ] = 8'h00;
    rom[ 869 ] = 8'h00;
    rom[ 870 ] = 8'h01;
    rom[ 871 ] = 8'h01;
    rom[ 872 ] = 8'h01;
    rom[ 873 ] = 8'h01;
    rom[ 874 ] = 8'h05;
    rom[ 875 ] = 8'h07;
    rom[ 876 ] = 8'h07;
    rom[ 877 ] = 8'h37;
    rom[ 878 ] = 8'h3F;
    rom[ 879 ] = 8'h3F;
    rom[ 880 ] = 8'h3F;
    rom[ 881 ] = 8'h3F;
    rom[ 882 ] = 8'h3F;
    rom[ 883 ] = 8'h3F;
    rom[ 884 ] = 8'hBF;
    rom[ 885 ] = 8'hFF;
    rom[ 886 ] = 8'hFF;
    rom[ 887 ] = 8'hFF;
    rom[ 888 ] = 8'hFF;
    rom[ 889 ] = 8'hFF;
    rom[ 890 ] = 8'hFF;
    rom[ 891 ] = 8'hFF;
    rom[ 892 ] = 8'hFF;
    rom[ 893 ] = 8'hFF;
    rom[ 894 ] = 8'hFF;
    rom[ 895 ] = 8'hFF;
    rom[ 896 ] = 8'hFF;
    rom[ 897 ] = 8'hFF;
    rom[ 898 ] = 8'hFF;
    rom[ 899 ] = 8'hFF;
    rom[ 900 ] = 8'hFF;
    rom[ 901 ] = 8'hFF;
    rom[ 902 ] = 8'hFF;
    rom[ 903 ] = 8'hFF;
    rom[ 904 ] = 8'hFF;
    rom[ 905 ] = 8'hFF;
    rom[ 906 ] = 8'hFF;
    rom[ 907 ] = 8'hFF;
    rom[ 908 ] = 8'hFF;
    rom[ 909 ] = 8'hFF;
    rom[ 910 ] = 8'hFF;
    rom[ 911 ] = 8'hFF;
    rom[ 912 ] = 8'hFF;
    rom[ 913 ] = 8'hFF;
    rom[ 914 ] = 8'hFF;
    rom[ 915 ] = 8'hFF;
    rom[ 916 ] = 8'hFF;
    rom[ 917 ] = 8'hFF;
    rom[ 918 ] = 8'hFF;
    rom[ 919 ] = 8'hFF;
    rom[ 920 ] = 8'hFF;
    rom[ 921 ] = 8'hFF;
    rom[ 922 ] = 8'hFF;
    rom[ 923 ] = 8'h3F;
    rom[ 924 ] = 8'h3F;
    rom[ 925 ] = 8'h3F;
    rom[ 926 ] = 8'h3F;
    rom[ 927 ] = 8'h3F;
    rom[ 928 ] = 8'h3F;
    rom[ 929 ] = 8'h3F;
    rom[ 930 ] = 8'h3F;
    rom[ 931 ] = 8'h3F;
    rom[ 932 ] = 8'h3F;
    rom[ 933 ] = 8'h3F;
    rom[ 934 ] = 8'h3F;
    rom[ 935 ] = 8'h3F;
    rom[ 936 ] = 8'h3F;
    rom[ 937 ] = 8'h3F;
    rom[ 938 ] = 8'h3F;
    rom[ 939 ] = 8'h3F;
    rom[ 940 ] = 8'h3F;
    rom[ 941 ] = 8'h3F;
    rom[ 942 ] = 8'h3F;
    rom[ 943 ] = 8'hFF;
    rom[ 944 ] = 8'hFF;
    rom[ 945 ] = 8'hFF;
    rom[ 946 ] = 8'hFF;
    rom[ 947 ] = 8'hFF;
    rom[ 948 ] = 8'hFF;
    rom[ 949 ] = 8'hFF;
    rom[ 950 ] = 8'hFF;
    rom[ 951 ] = 8'hFF;
    rom[ 952 ] = 8'hFF;
    rom[ 953 ] = 8'hFF;
    rom[ 954 ] = 8'hFF;
    rom[ 955 ] = 8'hFF;
    rom[ 956 ] = 8'hFF;
    rom[ 957 ] = 8'hFF;
    rom[ 958 ] = 8'hFF;
    rom[ 959 ] = 8'hFF;
    rom[ 960 ] = 8'hFF;
    rom[ 961 ] = 8'hFF;
    rom[ 962 ] = 8'hFF;
    rom[ 963 ] = 8'hFF;
    rom[ 964 ] = 8'hFF;
    rom[ 965 ] = 8'hFF;
    rom[ 966 ] = 8'hFF;
    rom[ 967 ] = 8'hFF;
    rom[ 968 ] = 8'hFF;
    rom[ 969 ] = 8'hFF;
    rom[ 970 ] = 8'hFF;
    rom[ 971 ] = 8'hFF;
    rom[ 972 ] = 8'hFF;
    rom[ 973 ] = 8'hFF;
    rom[ 974 ] = 8'hFF;
    rom[ 975 ] = 8'hFF;
    rom[ 976 ] = 8'hFF;
    rom[ 977 ] = 8'hFF;
    rom[ 978 ] = 8'hFF;
    rom[ 979 ] = 8'hFF;
    rom[ 980 ] = 8'hFF;
    rom[ 981 ] = 8'h7F;
    rom[ 982 ] = 8'h3F;
    rom[ 983 ] = 8'h3F;
    rom[ 984 ] = 8'h3F;
    rom[ 985 ] = 8'h3F;
    rom[ 986 ] = 8'h3F;
    rom[ 987 ] = 8'h3F;
    rom[ 988 ] = 8'h3F;
    rom[ 989 ] = 8'h3F;
    rom[ 990 ] = 8'h3F;
    rom[ 991 ] = 8'h3F;
    rom[ 992 ] = 8'h3F;
    rom[ 993 ] = 8'h3F;
    rom[ 994 ] = 8'h3F;
    rom[ 995 ] = 8'h3F;
    rom[ 996 ] = 8'h3F;
    rom[ 997 ] = 8'h3F;
    rom[ 998 ] = 8'h3F;
    rom[ 999 ] = 8'h3F;
    rom[1000 ] = 8'h3F;
    rom[1001 ] = 8'h3F;
    rom[1002 ] = 8'h3F;
    rom[1003 ] = 8'h3F;
    rom[1004 ] = 8'h3F;
    rom[1005 ] = 8'h3F;
    rom[1006 ] = 8'h3F;
    rom[1007 ] = 8'h3F;
    rom[1008 ] = 8'h3F;
    rom[1009 ] = 8'h3F;
    rom[1010 ] = 8'h3F;
    rom[1011 ] = 8'h3F;
    rom[1012 ] = 8'h3F;
    rom[1013 ] = 8'h3F;
    rom[1014 ] = 8'h0F;
    rom[1015 ] = 8'h03;
    rom[1016 ] = 8'h00;
    rom[1017 ] = 8'h00;
    rom[1018 ] = 8'h00;
    rom[1019 ] = 8'h00;
    rom[1020 ] = 8'h00;
    rom[1021 ] = 8'h00;
    rom[1022 ] = 8'h00;
    rom[1023 ] = 8'h00;
    rom[1024 ] = 8'h00;
    rom[1025 ] = 8'h00;
    rom[1026 ] = 8'h00;
    rom[1027 ] = 8'h00;
    rom[1028 ] = 8'h00;
    rom[1029 ] = 8'h00;
    rom[1030 ] = 8'h00;
    rom[1031 ] = 8'h00;
    rom[1032 ] = 8'h00;
    rom[1033 ] = 8'h00;
    rom[1034 ] = 8'h00;
    rom[1035 ] = 8'h00;
    rom[1036 ] = 8'h00;
    rom[1037 ] = 8'h00;
    rom[1038 ] = 8'h00;
    rom[1039 ] = 8'h00;
    rom[1040 ] = 8'h00;
    rom[1041 ] = 8'h00;
    rom[1042 ] = 8'h00;
    rom[1043 ] = 8'h00;
    rom[1044 ] = 8'h00;
    rom[1045 ] = 8'h00;
    rom[1046 ] = 8'h00;
    rom[1047 ] = 8'h00;
    rom[1048 ] = 8'h00;
    rom[1049 ] = 8'h00;
    rom[1050 ] = 8'h00;
    rom[1051 ] = 8'h00;
    rom[1052 ] = 8'h00;
    rom[1053 ] = 8'h00;
    rom[1054 ] = 8'h00;
    rom[1055 ] = 8'h00;
    rom[1056 ] = 8'h00;
    rom[1057 ] = 8'h00;
    rom[1058 ] = 8'h00;
    rom[1059 ] = 8'h00;
    rom[1060 ] = 8'h00;
    rom[1061 ] = 8'h00;
    rom[1062 ] = 8'h00;
    rom[1063 ] = 8'h00;
    rom[1064 ] = 8'h00;
    rom[1065 ] = 8'h00;
    rom[1066 ] = 8'h00;
    rom[1067 ] = 8'h00;
    rom[1068 ] = 8'h00;
    rom[1069 ] = 8'hC0;
    rom[1070 ] = 8'hF0;
    rom[1071 ] = 8'hFC;
    rom[1072 ] = 8'hFE;
    rom[1073 ] = 8'hFE;
    rom[1074 ] = 8'hFE;
    rom[1075 ] = 8'hFE;
    rom[1076 ] = 8'hFE;
    rom[1077 ] = 8'hFE;
    rom[1078 ] = 8'hFE;
    rom[1079 ] = 8'hFE;
    rom[1080 ] = 8'hFE;
    rom[1081 ] = 8'hFE;
    rom[1082 ] = 8'hFE;
    rom[1083 ] = 8'hFE;
    rom[1084 ] = 8'hFE;
    rom[1085 ] = 8'hFE;
    rom[1086 ] = 8'hFE;
    rom[1087 ] = 8'hFE;
    rom[1088 ] = 8'hFE;
    rom[1089 ] = 8'hFE;
    rom[1090 ] = 8'hFE;
    rom[1091 ] = 8'hFE;
    rom[1092 ] = 8'hFE;
    rom[1093 ] = 8'hFE;
    rom[1094 ] = 8'hFE;
    rom[1095 ] = 8'hFE;
    rom[1096 ] = 8'hFE;
    rom[1097 ] = 8'hFE;
    rom[1098 ] = 8'hFE;
    rom[1099 ] = 8'hFE;
    rom[1100 ] = 8'hF0;
    rom[1101 ] = 8'hF0;
    rom[1102 ] = 8'hF0;
    rom[1103 ] = 8'hC0;
    rom[1104 ] = 8'hC0;
    rom[1105 ] = 8'hC0;
    rom[1106 ] = 8'hC0;
    rom[1107 ] = 8'h40;
    rom[1108 ] = 8'h00;
    rom[1109 ] = 8'h00;
    rom[1110 ] = 8'h00;
    rom[1111 ] = 8'h00;
    rom[1112 ] = 8'h00;
    rom[1113 ] = 8'h00;
    rom[1114 ] = 8'h00;
    rom[1115 ] = 8'h00;
    rom[1116 ] = 8'h00;
    rom[1117 ] = 8'h00;
    rom[1118 ] = 8'h00;
    rom[1119 ] = 8'h00;
    rom[1120 ] = 8'h00;
    rom[1121 ] = 8'h00;
    rom[1122 ] = 8'h00;
    rom[1123 ] = 8'h00;
    rom[1124 ] = 8'h00;
    rom[1125 ] = 8'h00;
    rom[1126 ] = 8'h00;
    rom[1127 ] = 8'h00;
    rom[1128 ] = 8'h00;
    rom[1129 ] = 8'h00;
    rom[1130 ] = 8'h00;
    rom[1131 ] = 8'h00;
    rom[1132 ] = 8'h00;
    rom[1133 ] = 8'h00;
    rom[1134 ] = 8'h80;
    rom[1135 ] = 8'hC0;
    rom[1136 ] = 8'hC0;
    rom[1137 ] = 8'hF0;
    rom[1138 ] = 8'hFC;
    rom[1139 ] = 8'hFF;
    rom[1140 ] = 8'hFF;
    rom[1141 ] = 8'hFF;
    rom[1142 ] = 8'hFF;
    rom[1143 ] = 8'hFF;
    rom[1144 ] = 8'hFF;
    rom[1145 ] = 8'hFF;
    rom[1146 ] = 8'hFF;
    rom[1147 ] = 8'hFF;
    rom[1148 ] = 8'hFF;
    rom[1149 ] = 8'hFF;
    rom[1150 ] = 8'hFF;
    rom[1151 ] = 8'hFF;
    rom[1152 ] = 8'hFF;
    rom[1153 ] = 8'hFF;
    rom[1154 ] = 8'hFF;
    rom[1155 ] = 8'hFF;
    rom[1156 ] = 8'hFF;
    rom[1157 ] = 8'hFF;
    rom[1158 ] = 8'hFF;
    rom[1159 ] = 8'hFF;
    rom[1160 ] = 8'hFF;
    rom[1161 ] = 8'hFF;
    rom[1162 ] = 8'hFF;
    rom[1163 ] = 8'hFF;
    rom[1164 ] = 8'hFF;
    rom[1165 ] = 8'hFF;
    rom[1166 ] = 8'hFF;
    rom[1167 ] = 8'hFF;
    rom[1168 ] = 8'hFF;
    rom[1169 ] = 8'hFF;
    rom[1170 ] = 8'hFF;
    rom[1171 ] = 8'hFF;
    rom[1172 ] = 8'hFF;
    rom[1173 ] = 8'hFF;
    rom[1174 ] = 8'h7F;
    rom[1175 ] = 8'h1F;
    rom[1176 ] = 8'h0F;
    rom[1177 ] = 8'h03;
    rom[1178 ] = 8'h00;
    rom[1179 ] = 8'h00;
    rom[1180 ] = 8'h00;
    rom[1181 ] = 8'h00;
    rom[1182 ] = 8'h00;
    rom[1183 ] = 8'h00;
    rom[1184 ] = 8'h00;
    rom[1185 ] = 8'h00;
    rom[1186 ] = 8'h00;
    rom[1187 ] = 8'h00;
    rom[1188 ] = 8'h00;
    rom[1189 ] = 8'h00;
    rom[1190 ] = 8'h00;
    rom[1191 ] = 8'h00;
    rom[1192 ] = 8'h00;
    rom[1193 ] = 8'h00;
    rom[1194 ] = 8'h80;
    rom[1195 ] = 8'hE0;
    rom[1196 ] = 8'hF8;
    rom[1197 ] = 8'hFC;
    rom[1198 ] = 8'hFF;
    rom[1199 ] = 8'hFF;
    rom[1200 ] = 8'hFF;
    rom[1201 ] = 8'hFF;
    rom[1202 ] = 8'hFF;
    rom[1203 ] = 8'hFF;
    rom[1204 ] = 8'hFF;
    rom[1205 ] = 8'hFF;
    rom[1206 ] = 8'hFF;
    rom[1207 ] = 8'hFF;
    rom[1208 ] = 8'hFF;
    rom[1209 ] = 8'hFF;
    rom[1210 ] = 8'hFF;
    rom[1211 ] = 8'hFF;
    rom[1212 ] = 8'hFF;
    rom[1213 ] = 8'hFF;
    rom[1214 ] = 8'hFF;
    rom[1215 ] = 8'hFF;
    rom[1216 ] = 8'hFF;
    rom[1217 ] = 8'hFF;
    rom[1218 ] = 8'hFF;
    rom[1219 ] = 8'hFF;
    rom[1220 ] = 8'hFF;
    rom[1221 ] = 8'hFF;
    rom[1222 ] = 8'hFF;
    rom[1223 ] = 8'hFF;
    rom[1224 ] = 8'hFF;
    rom[1225 ] = 8'hFF;
    rom[1226 ] = 8'hFF;
    rom[1227 ] = 8'hFF;
    rom[1228 ] = 8'hFF;
    rom[1229 ] = 8'hFF;
    rom[1230 ] = 8'hFF;
    rom[1231 ] = 8'hFF;
    rom[1232 ] = 8'hFF;
    rom[1233 ] = 8'h7F;
    rom[1234 ] = 8'h1F;
    rom[1235 ] = 8'h07;
    rom[1236 ] = 8'h01;
    rom[1237 ] = 8'h00;
    rom[1238 ] = 8'h00;
    rom[1239 ] = 8'h00;
    rom[1240 ] = 8'h00;
    rom[1241 ] = 8'h00;
    rom[1242 ] = 8'h00;
    rom[1243 ] = 8'h00;
    rom[1244 ] = 8'h00;
    rom[1245 ] = 8'h00;
    rom[1246 ] = 8'h00;
    rom[1247 ] = 8'h00;
    rom[1248 ] = 8'h00;
    rom[1249 ] = 8'h00;
    rom[1250 ] = 8'h00;
    rom[1251 ] = 8'h00;
    rom[1252 ] = 8'h00;
    rom[1253 ] = 8'h00;
    rom[1254 ] = 8'h00;
    rom[1255 ] = 8'h00;
    rom[1256 ] = 8'h00;
    rom[1257 ] = 8'h00;
    rom[1258 ] = 8'h00;
    rom[1259 ] = 8'h00;
    rom[1260 ] = 8'h00;
    rom[1261 ] = 8'h00;
    rom[1262 ] = 8'h00;
    rom[1263 ] = 8'h00;
    rom[1264 ] = 8'h00;
    rom[1265 ] = 8'h00;
    rom[1266 ] = 8'h00;
    rom[1267 ] = 8'h00;
    rom[1268 ] = 8'h00;
    rom[1269 ] = 8'h00;
    rom[1270 ] = 8'h00;
    rom[1271 ] = 8'h00;
    rom[1272 ] = 8'h00;
    rom[1273 ] = 8'h00;
    rom[1274 ] = 8'h00;
    rom[1275 ] = 8'h00;
    rom[1276 ] = 8'h00;
    rom[1277 ] = 8'h00;
    rom[1278 ] = 8'h00;
    rom[1279 ] = 8'h00;
    rom[1280 ] = 8'h00;
    rom[1281 ] = 8'h00;
    rom[1282 ] = 8'h00;
    rom[1283 ] = 8'h00;
    rom[1284 ] = 8'h00;
    rom[1285 ] = 8'h00;
    rom[1286 ] = 8'h00;
    rom[1287 ] = 8'h00;
    rom[1288 ] = 8'h00;
    rom[1289 ] = 8'h00;
    rom[1290 ] = 8'h00;
    rom[1291 ] = 8'h00;
    rom[1292 ] = 8'h00;
    rom[1293 ] = 8'h00;
    rom[1294 ] = 8'h00;
    rom[1295 ] = 8'h00;
    rom[1296 ] = 8'h00;
    rom[1297 ] = 8'h00;
    rom[1298 ] = 8'h00;
    rom[1299 ] = 8'h00;
    rom[1300 ] = 8'h00;
    rom[1301 ] = 8'h00;
    rom[1302 ] = 8'h00;
    rom[1303 ] = 8'h00;
    rom[1304 ] = 8'h00;
    rom[1305 ] = 8'h00;
    rom[1306 ] = 8'h00;
    rom[1307 ] = 8'h00;
    rom[1308 ] = 8'h00;
    rom[1309 ] = 8'h00;
    rom[1310 ] = 8'h00;
    rom[1311 ] = 8'h00;
    rom[1312 ] = 8'h00;
    rom[1313 ] = 8'h00;
    rom[1314 ] = 8'h00;
    rom[1315 ] = 8'h00;
    rom[1316 ] = 8'h00;
    rom[1317 ] = 8'h00;
    rom[1318 ] = 8'h00;
    rom[1319 ] = 8'h00;
    rom[1320 ] = 8'h00;
    rom[1321 ] = 8'h00;
    rom[1322 ] = 8'h00;
    rom[1323 ] = 8'h00;
    rom[1324 ] = 8'h00;
    rom[1325 ] = 8'h3F;
    rom[1326 ] = 8'h7F;
    rom[1327 ] = 8'hFF;
    rom[1328 ] = 8'hFF;
    rom[1329 ] = 8'hFF;
    rom[1330 ] = 8'hFF;
    rom[1331 ] = 8'hFF;
    rom[1332 ] = 8'hFF;
    rom[1333 ] = 8'hFF;
    rom[1334 ] = 8'hFF;
    rom[1335 ] = 8'hFF;
    rom[1336 ] = 8'hFF;
    rom[1337 ] = 8'hFF;
    rom[1338 ] = 8'hFF;
    rom[1339 ] = 8'hFF;
    rom[1340 ] = 8'hFF;
    rom[1341 ] = 8'hFF;
    rom[1342 ] = 8'hFF;
    rom[1343 ] = 8'hFF;
    rom[1344 ] = 8'hFF;
    rom[1345 ] = 8'hFF;
    rom[1346 ] = 8'hFF;
    rom[1347 ] = 8'hFF;
    rom[1348 ] = 8'hFF;
    rom[1349 ] = 8'hFF;
    rom[1350 ] = 8'hFF;
    rom[1351 ] = 8'hFF;
    rom[1352 ] = 8'hFF;
    rom[1353 ] = 8'hFF;
    rom[1354 ] = 8'hFF;
    rom[1355 ] = 8'hFF;
    rom[1356 ] = 8'hFF;
    rom[1357 ] = 8'hFF;
    rom[1358 ] = 8'hFF;
    rom[1359 ] = 8'hFF;
    rom[1360 ] = 8'hFF;
    rom[1361 ] = 8'hFF;
    rom[1362 ] = 8'hF9;
    rom[1363 ] = 8'hF8;
    rom[1364 ] = 8'hF8;
    rom[1365 ] = 8'hF8;
    rom[1366 ] = 8'hF8;
    rom[1367 ] = 8'hF8;
    rom[1368 ] = 8'hF8;
    rom[1369 ] = 8'hF8;
    rom[1370 ] = 8'hF8;
    rom[1371 ] = 8'hF8;
    rom[1372 ] = 8'hF8;
    rom[1373 ] = 8'hF8;
    rom[1374 ] = 8'hF8;
    rom[1375 ] = 8'hF8;
    rom[1376 ] = 8'hF8;
    rom[1377 ] = 8'hF8;
    rom[1378 ] = 8'hF8;
    rom[1379 ] = 8'hF8;
    rom[1380 ] = 8'hFC;
    rom[1381 ] = 8'hFC;
    rom[1382 ] = 8'hFC;
    rom[1383 ] = 8'hFC;
    rom[1384 ] = 8'hFC;
    rom[1385 ] = 8'hFE;
    rom[1386 ] = 8'hFE;
    rom[1387 ] = 8'hFE;
    rom[1388 ] = 8'hFF;
    rom[1389 ] = 8'hFF;
    rom[1390 ] = 8'hFF;
    rom[1391 ] = 8'hFF;
    rom[1392 ] = 8'hFF;
    rom[1393 ] = 8'hFF;
    rom[1394 ] = 8'hFF;
    rom[1395 ] = 8'hFF;
    rom[1396 ] = 8'hFF;
    rom[1397 ] = 8'hFF;
    rom[1398 ] = 8'hFF;
    rom[1399 ] = 8'hFF;
    rom[1400 ] = 8'hFF;
    rom[1401 ] = 8'hFF;
    rom[1402 ] = 8'hFF;
    rom[1403 ] = 8'hFF;
    rom[1404 ] = 8'hFF;
    rom[1405 ] = 8'hFF;
    rom[1406 ] = 8'hFF;
    rom[1407 ] = 8'hFF;
    rom[1408 ] = 8'hFF;
    rom[1409 ] = 8'hFF;
    rom[1410 ] = 8'hFF;
    rom[1411 ] = 8'hFF;
    rom[1412 ] = 8'hFF;
    rom[1413 ] = 8'hFF;
    rom[1414 ] = 8'hFF;
    rom[1415 ] = 8'hFF;
    rom[1416 ] = 8'hFF;
    rom[1417 ] = 8'hFF;
    rom[1418 ] = 8'hFF;
    rom[1419 ] = 8'hFF;
    rom[1420 ] = 8'hFF;
    rom[1421 ] = 8'hFF;
    rom[1422 ] = 8'hFF;
    rom[1423 ] = 8'hFF;
    rom[1424 ] = 8'hFF;
    rom[1425 ] = 8'h7F;
    rom[1426 ] = 8'h3F;
    rom[1427 ] = 8'h1F;
    rom[1428 ] = 8'h07;
    rom[1429 ] = 8'h01;
    rom[1430 ] = 8'h00;
    rom[1431 ] = 8'h00;
    rom[1432 ] = 8'h00;
    rom[1433 ] = 8'h00;
    rom[1434 ] = 8'h00;
    rom[1435 ] = 8'h00;
    rom[1436 ] = 8'h00;
    rom[1437 ] = 8'h00;
    rom[1438 ] = 8'h00;
    rom[1439 ] = 8'h00;
    rom[1440 ] = 8'h00;
    rom[1441 ] = 8'h00;
    rom[1442 ] = 8'h00;
    rom[1443 ] = 8'h00;
    rom[1444 ] = 8'h00;
    rom[1445 ] = 8'h00;
    rom[1446 ] = 8'h80;
    rom[1447 ] = 8'hE0;
    rom[1448 ] = 8'hF8;
    rom[1449 ] = 8'hFE;
    rom[1450 ] = 8'hFF;
    rom[1451 ] = 8'hFF;
    rom[1452 ] = 8'hFF;
    rom[1453 ] = 8'hFF;
    rom[1454 ] = 8'hFF;
    rom[1455 ] = 8'hFF;
    rom[1456 ] = 8'hFF;
    rom[1457 ] = 8'hFF;
    rom[1458 ] = 8'hFF;
    rom[1459 ] = 8'hFF;
    rom[1460 ] = 8'hFF;
    rom[1461 ] = 8'hFF;
    rom[1462 ] = 8'hFF;
    rom[1463 ] = 8'hFF;
    rom[1464 ] = 8'hFF;
    rom[1465 ] = 8'hFF;
    rom[1466 ] = 8'hFF;
    rom[1467 ] = 8'hFF;
    rom[1468 ] = 8'hFF;
    rom[1469 ] = 8'hFF;
    rom[1470 ] = 8'hFF;
    rom[1471 ] = 8'hFF;
    rom[1472 ] = 8'hFF;
    rom[1473 ] = 8'hFF;
    rom[1474 ] = 8'hFF;
    rom[1475 ] = 8'hFF;
    rom[1476 ] = 8'hFF;
    rom[1477 ] = 8'hFF;
    rom[1478 ] = 8'hFF;
    rom[1479 ] = 8'hFF;
    rom[1480 ] = 8'hFF;
    rom[1481 ] = 8'hFF;
    rom[1482 ] = 8'hFF;
    rom[1483 ] = 8'hFF;
    rom[1484 ] = 8'hFF;
    rom[1485 ] = 8'h3F;
    rom[1486 ] = 8'h0F;
    rom[1487 ] = 8'h03;
    rom[1488 ] = 8'h00;
    rom[1489 ] = 8'h00;
    rom[1490 ] = 8'h00;
    rom[1491 ] = 8'h00;
    rom[1492 ] = 8'h00;
    rom[1493 ] = 8'h00;
    rom[1494 ] = 8'h00;
    rom[1495 ] = 8'h00;
    rom[1496 ] = 8'h00;
    rom[1497 ] = 8'h00;
    rom[1498 ] = 8'h00;
    rom[1499 ] = 8'h00;
    rom[1500 ] = 8'h00;
    rom[1501 ] = 8'h00;
    rom[1502 ] = 8'h00;
    rom[1503 ] = 8'h00;
    rom[1504 ] = 8'h00;
    rom[1505 ] = 8'h00;
    rom[1506 ] = 8'h00;
    rom[1507 ] = 8'h00;
    rom[1508 ] = 8'h00;
    rom[1509 ] = 8'h00;
    rom[1510 ] = 8'h00;
    rom[1511 ] = 8'h00;
    rom[1512 ] = 8'h00;
    rom[1513 ] = 8'h00;
    rom[1514 ] = 8'h00;
    rom[1515 ] = 8'h00;
    rom[1516 ] = 8'h00;
    rom[1517 ] = 8'h00;
    rom[1518 ] = 8'h00;
    rom[1519 ] = 8'h00;
    rom[1520 ] = 8'h00;
    rom[1521 ] = 8'h00;
    rom[1522 ] = 8'h00;
    rom[1523 ] = 8'h00;
    rom[1524 ] = 8'h00;
    rom[1525 ] = 8'h00;
    rom[1526 ] = 8'h00;
    rom[1527 ] = 8'h00;
    rom[1528 ] = 8'h00;
    rom[1529 ] = 8'h00;
    rom[1530 ] = 8'h00;
    rom[1531 ] = 8'h00;
    rom[1532 ] = 8'h00;
    rom[1533 ] = 8'h00;
    rom[1534 ] = 8'h00;
    rom[1535 ] = 8'h00;
    rom[1536 ] = 8'h00;
    rom[1537 ] = 8'h00;
    rom[1538 ] = 8'h00;
    rom[1539 ] = 8'h00;
    rom[1540 ] = 8'h00;
    rom[1541 ] = 8'h00;
    rom[1542 ] = 8'h00;
    rom[1543 ] = 8'h00;
    rom[1544 ] = 8'h00;
    rom[1545 ] = 8'h00;
    rom[1546 ] = 8'h00;
    rom[1547 ] = 8'h00;
    rom[1548 ] = 8'h00;
    rom[1549 ] = 8'h00;
    rom[1550 ] = 8'h00;
    rom[1551 ] = 8'h00;
    rom[1552 ] = 8'h00;
    rom[1553 ] = 8'h00;
    rom[1554 ] = 8'h00;
    rom[1555 ] = 8'h00;
    rom[1556 ] = 8'h00;
    rom[1557 ] = 8'h00;
    rom[1558 ] = 8'h00;
    rom[1559 ] = 8'h00;
    rom[1560 ] = 8'h00;
    rom[1561 ] = 8'h00;
    rom[1562 ] = 8'h00;
    rom[1563 ] = 8'h00;
    rom[1564 ] = 8'h00;
    rom[1565 ] = 8'h00;
    rom[1566 ] = 8'h00;
    rom[1567 ] = 8'h00;
    rom[1568 ] = 8'h00;
    rom[1569 ] = 8'h00;
    rom[1570 ] = 8'h00;
    rom[1571 ] = 8'h00;
    rom[1572 ] = 8'h00;
    rom[1573 ] = 8'h00;
    rom[1574 ] = 8'h00;
    rom[1575 ] = 8'h00;
    rom[1576 ] = 8'h00;
    rom[1577 ] = 8'h00;
    rom[1578 ] = 8'h00;
    rom[1579 ] = 8'h00;
    rom[1580 ] = 8'h00;
    rom[1581 ] = 8'h00;
    rom[1582 ] = 8'h00;
    rom[1583 ] = 8'h01;
    rom[1584 ] = 8'h03;
    rom[1585 ] = 8'h03;
    rom[1586 ] = 8'h07;
    rom[1587 ] = 8'h0F;
    rom[1588 ] = 8'h0F;
    rom[1589 ] = 8'h1F;
    rom[1590 ] = 8'h1F;
    rom[1591 ] = 8'h3F;
    rom[1592 ] = 8'h3F;
    rom[1593 ] = 8'h7F;
    rom[1594 ] = 8'hFF;
    rom[1595 ] = 8'hFF;
    rom[1596 ] = 8'hFF;
    rom[1597 ] = 8'hFF;
    rom[1598 ] = 8'hFF;
    rom[1599 ] = 8'hFF;
    rom[1600 ] = 8'hFF;
    rom[1601 ] = 8'hFF;
    rom[1602 ] = 8'hFF;
    rom[1603 ] = 8'hFF;
    rom[1604 ] = 8'hFF;
    rom[1605 ] = 8'hFF;
    rom[1606 ] = 8'hFF;
    rom[1607 ] = 8'hFF;
    rom[1608 ] = 8'hFF;
    rom[1609 ] = 8'hFF;
    rom[1610 ] = 8'hFF;
    rom[1611 ] = 8'hFF;
    rom[1612 ] = 8'hFF;
    rom[1613 ] = 8'hFF;
    rom[1614 ] = 8'hFF;
    rom[1615 ] = 8'hFF;
    rom[1616 ] = 8'hFF;
    rom[1617 ] = 8'hFF;
    rom[1618 ] = 8'hFF;
    rom[1619 ] = 8'hFF;
    rom[1620 ] = 8'hFF;
    rom[1621 ] = 8'hFF;
    rom[1622 ] = 8'hFF;
    rom[1623 ] = 8'hFF;
    rom[1624 ] = 8'hFF;
    rom[1625 ] = 8'hFF;
    rom[1626 ] = 8'hFF;
    rom[1627 ] = 8'hFF;
    rom[1628 ] = 8'hFF;
    rom[1629 ] = 8'hFF;
    rom[1630 ] = 8'hFF;
    rom[1631 ] = 8'hFF;
    rom[1632 ] = 8'hFF;
    rom[1633 ] = 8'hFF;
    rom[1634 ] = 8'hFF;
    rom[1635 ] = 8'hFF;
    rom[1636 ] = 8'hFF;
    rom[1637 ] = 8'hFF;
    rom[1638 ] = 8'hFF;
    rom[1639 ] = 8'hFF;
    rom[1640 ] = 8'hFF;
    rom[1641 ] = 8'hFF;
    rom[1642 ] = 8'hFF;
    rom[1643 ] = 8'hFF;
    rom[1644 ] = 8'hFF;
    rom[1645 ] = 8'hFF;
    rom[1646 ] = 8'hFF;
    rom[1647 ] = 8'hFF;
    rom[1648 ] = 8'hFF;
    rom[1649 ] = 8'hFF;
    rom[1650 ] = 8'hFF;
    rom[1651 ] = 8'hFF;
    rom[1652 ] = 8'hFF;
    rom[1653 ] = 8'hFF;
    rom[1654 ] = 8'hFF;
    rom[1655 ] = 8'hFF;
    rom[1656 ] = 8'hFF;
    rom[1657 ] = 8'hFF;
    rom[1658 ] = 8'hFF;
    rom[1659 ] = 8'hFF;
    rom[1660 ] = 8'hFF;
    rom[1661 ] = 8'hFF;
    rom[1662 ] = 8'hFF;
    rom[1663 ] = 8'hFF;
    rom[1664 ] = 8'hFF;
    rom[1665 ] = 8'hFF;
    rom[1666 ] = 8'hFF;
    rom[1667 ] = 8'hFF;
    rom[1668 ] = 8'h7F;
    rom[1669 ] = 8'h7F;
    rom[1670 ] = 8'h3F;
    rom[1671 ] = 8'h3F;
    rom[1672 ] = 8'h1F;
    rom[1673 ] = 8'h1F;
    rom[1674 ] = 8'h0F;
    rom[1675 ] = 8'h0F;
    rom[1676 ] = 8'h07;
    rom[1677 ] = 8'h03;
    rom[1678 ] = 8'h03;
    rom[1679 ] = 8'h01;
    rom[1680 ] = 8'h00;
    rom[1681 ] = 8'h00;
    rom[1682 ] = 8'h00;
    rom[1683 ] = 8'h00;
    rom[1684 ] = 8'h00;
    rom[1685 ] = 8'h00;
    rom[1686 ] = 8'h00;
    rom[1687 ] = 8'h00;
    rom[1688 ] = 8'h00;
    rom[1689 ] = 8'h00;
    rom[1690 ] = 8'h00;
    rom[1691 ] = 8'h00;
    rom[1692 ] = 8'h00;
    rom[1693 ] = 8'h00;
    rom[1694 ] = 8'h00;
    rom[1695 ] = 8'h00;
    rom[1696 ] = 8'h00;
    rom[1697 ] = 8'h00;
    rom[1698 ] = 8'hC0;
    rom[1699 ] = 8'hF0;
    rom[1700 ] = 8'hFC;
    rom[1701 ] = 8'hFF;
    rom[1702 ] = 8'hFF;
    rom[1703 ] = 8'hFF;
    rom[1704 ] = 8'hFF;
    rom[1705 ] = 8'hFF;
    rom[1706 ] = 8'hFF;
    rom[1707 ] = 8'hFF;
    rom[1708 ] = 8'hFF;
    rom[1709 ] = 8'hFF;
    rom[1710 ] = 8'hFF;
    rom[1711 ] = 8'hFF;
    rom[1712 ] = 8'hFF;
    rom[1713 ] = 8'hFF;
    rom[1714 ] = 8'hFF;
    rom[1715 ] = 8'hFF;
    rom[1716 ] = 8'hFF;
    rom[1717 ] = 8'hFF;
    rom[1718 ] = 8'hFF;
    rom[1719 ] = 8'hFF;
    rom[1720 ] = 8'hFF;
    rom[1721 ] = 8'hFF;
    rom[1722 ] = 8'hFF;
    rom[1723 ] = 8'hFF;
    rom[1724 ] = 8'hFF;
    rom[1725 ] = 8'hFF;
    rom[1726 ] = 8'hFF;
    rom[1727 ] = 8'hFF;
    rom[1728 ] = 8'hFF;
    rom[1729 ] = 8'hFF;
    rom[1730 ] = 8'hFF;
    rom[1731 ] = 8'hFF;
    rom[1732 ] = 8'hFF;
    rom[1733 ] = 8'hFF;
    rom[1734 ] = 8'hFF;
    rom[1735 ] = 8'hFF;
    rom[1736 ] = 8'h7F;
    rom[1737 ] = 8'h1F;
    rom[1738 ] = 8'h0F;
    rom[1739 ] = 8'h03;
    rom[1740 ] = 8'h00;
    rom[1741 ] = 8'h00;
    rom[1742 ] = 8'h00;
    rom[1743 ] = 8'h00;
    rom[1744 ] = 8'h00;
    rom[1745 ] = 8'h00;
    rom[1746 ] = 8'h00;
    rom[1747 ] = 8'h00;
    rom[1748 ] = 8'h00;
    rom[1749 ] = 8'h00;
    rom[1750 ] = 8'h00;
    rom[1751 ] = 8'h00;
    rom[1752 ] = 8'h00;
    rom[1753 ] = 8'h00;
    rom[1754 ] = 8'h00;
    rom[1755 ] = 8'h00;
    rom[1756 ] = 8'h00;
    rom[1757 ] = 8'h00;
    rom[1758 ] = 8'h00;
    rom[1759 ] = 8'h00;
    rom[1760 ] = 8'h00;
    rom[1761 ] = 8'h00;
    rom[1762 ] = 8'h00;
    rom[1763 ] = 8'h00;
    rom[1764 ] = 8'h00;
    rom[1765 ] = 8'h00;
    rom[1766 ] = 8'h00;
    rom[1767 ] = 8'h00;
    rom[1768 ] = 8'h00;
    rom[1769 ] = 8'h00;
    rom[1770 ] = 8'h00;
    rom[1771 ] = 8'h00;
    rom[1772 ] = 8'h00;
    rom[1773 ] = 8'h00;
    rom[1774 ] = 8'h00;
    rom[1775 ] = 8'h00;
    rom[1776 ] = 8'h00;
    rom[1777 ] = 8'h00;
    rom[1778 ] = 8'h00;
    rom[1779 ] = 8'h00;
    rom[1780 ] = 8'h00;
    rom[1781 ] = 8'h00;
    rom[1782 ] = 8'h00;
    rom[1783 ] = 8'h00;
    rom[1784 ] = 8'h00;
    rom[1785 ] = 8'h00;
    rom[1786 ] = 8'h00;
    rom[1787 ] = 8'h00;
    rom[1788 ] = 8'h00;
    rom[1789 ] = 8'h00;
    rom[1790 ] = 8'h00;
    rom[1791 ] = 8'h00;
    rom[1792 ] = 8'h00;
    rom[1793 ] = 8'h00;
    rom[1794 ] = 8'h00;
    rom[1795 ] = 8'h00;
    rom[1796 ] = 8'h00;
    rom[1797 ] = 8'h00;
    rom[1798 ] = 8'h00;
    rom[1799 ] = 8'h00;
    rom[1800 ] = 8'h00;
    rom[1801 ] = 8'h00;
    rom[1802 ] = 8'h00;
    rom[1803 ] = 8'h00;
    rom[1804 ] = 8'h00;
    rom[1805 ] = 8'h00;
    rom[1806 ] = 8'h00;
    rom[1807 ] = 8'h00;
    rom[1808 ] = 8'h00;
    rom[1809 ] = 8'h00;
    rom[1810 ] = 8'h00;
    rom[1811 ] = 8'h00;
    rom[1812 ] = 8'h00;
    rom[1813 ] = 8'h00;
    rom[1814 ] = 8'h00;
    rom[1815 ] = 8'h00;
    rom[1816 ] = 8'h00;
    rom[1817 ] = 8'h00;
    rom[1818 ] = 8'h00;
    rom[1819 ] = 8'h00;
    rom[1820 ] = 8'h00;
    rom[1821 ] = 8'h00;
    rom[1822 ] = 8'h00;
    rom[1823 ] = 8'h00;
    rom[1824 ] = 8'h00;
    rom[1825 ] = 8'h00;
    rom[1826 ] = 8'h00;
    rom[1827 ] = 8'h00;
    rom[1828 ] = 8'h00;
    rom[1829 ] = 8'h00;
    rom[1830 ] = 8'h00;
    rom[1831 ] = 8'h00;
    rom[1832 ] = 8'h00;
    rom[1833 ] = 8'h00;
    rom[1834 ] = 8'h00;
    rom[1835 ] = 8'h00;
    rom[1836 ] = 8'h00;
    rom[1837 ] = 8'h00;
    rom[1838 ] = 8'h00;
    rom[1839 ] = 8'h00;
    rom[1840 ] = 8'h00;
    rom[1841 ] = 8'h00;
    rom[1842 ] = 8'h00;
    rom[1843 ] = 8'h00;
    rom[1844 ] = 8'h00;
    rom[1845 ] = 8'h00;
    rom[1846 ] = 8'h00;
    rom[1847 ] = 8'h00;
    rom[1848 ] = 8'h00;
    rom[1849 ] = 8'h00;
    rom[1850 ] = 8'h00;
    rom[1851 ] = 8'h01;
    rom[1852 ] = 8'h01;
    rom[1853 ] = 8'h03;
    rom[1854 ] = 8'h03;
    rom[1855 ] = 8'h03;
    rom[1856 ] = 8'h07;
    rom[1857 ] = 8'h07;
    rom[1858 ] = 8'h07;
    rom[1859 ] = 8'h0F;
    rom[1860 ] = 8'h0F;
    rom[1861 ] = 8'h0F;
    rom[1862 ] = 8'h0F;
    rom[1863 ] = 8'h0F;
    rom[1864 ] = 8'h1F;
    rom[1865 ] = 8'h1F;
    rom[1866 ] = 8'h1F;
    rom[1867 ] = 8'h1F;
    rom[1868 ] = 8'h1F;
    rom[1869 ] = 8'h1F;
    rom[1870 ] = 8'h1F;
    rom[1871 ] = 8'h1F;
    rom[1872 ] = 8'h1F;
    rom[1873 ] = 8'h1F;
    rom[1874 ] = 8'h1F;
    rom[1875 ] = 8'h1F;
    rom[1876 ] = 8'h1F;
    rom[1877 ] = 8'h1F;
    rom[1878 ] = 8'h1F;
    rom[1879 ] = 8'h1F;
    rom[1880 ] = 8'h1F;
    rom[1881 ] = 8'h1F;
    rom[1882 ] = 8'h1F;
    rom[1883 ] = 8'h1F;
    rom[1884 ] = 8'h1F;
    rom[1885 ] = 8'h1F;
    rom[1886 ] = 8'h1F;
    rom[1887 ] = 8'h1F;
    rom[1888 ] = 8'h1F;
    rom[1889 ] = 8'h1F;
    rom[1890 ] = 8'h1F;
    rom[1891 ] = 8'h1F;
    rom[1892 ] = 8'h1F;
    rom[1893 ] = 8'h1F;
    rom[1894 ] = 8'h1F;
    rom[1895 ] = 8'h1F;
    rom[1896 ] = 8'h1F;
    rom[1897 ] = 8'h1F;
    rom[1898 ] = 8'h1F;
    rom[1899 ] = 8'h1F;
    rom[1900 ] = 8'h1F;
    rom[1901 ] = 8'h1F;
    rom[1902 ] = 8'h1F;
    rom[1903 ] = 8'h1F;
    rom[1904 ] = 8'h1F;
    rom[1905 ] = 8'h0F;
    rom[1906 ] = 8'h0F;
    rom[1907 ] = 8'h0F;
    rom[1908 ] = 8'h0F;
    rom[1909 ] = 8'h0F;
    rom[1910 ] = 8'h0F;
    rom[1911 ] = 8'h07;
    rom[1912 ] = 8'h07;
    rom[1913 ] = 8'h07;
    rom[1914 ] = 8'h07;
    rom[1915 ] = 8'h03;
    rom[1916 ] = 8'h03;
    rom[1917 ] = 8'h03;
    rom[1918 ] = 8'h01;
    rom[1919 ] = 8'h01;
    rom[1920 ] = 8'h01;
    rom[1921 ] = 8'h00;
    rom[1922 ] = 8'h00;
    rom[1923 ] = 8'h00;
    rom[1924 ] = 8'h00;
    rom[1925 ] = 8'h00;
    rom[1926 ] = 8'h00;
    rom[1927 ] = 8'h00;
    rom[1928 ] = 8'h00;
    rom[1929 ] = 8'h00;
    rom[1930 ] = 8'h00;
    rom[1931 ] = 8'h00;
    rom[1932 ] = 8'h00;
    rom[1933 ] = 8'h00;
    rom[1934 ] = 8'h00;
    rom[1935 ] = 8'h00;
    rom[1936 ] = 8'h00;
    rom[1937 ] = 8'h00;
    rom[1938 ] = 8'h00;
    rom[1939 ] = 8'h00;
    rom[1940 ] = 8'h00;
    rom[1941 ] = 8'h00;
    rom[1942 ] = 8'h00;
    rom[1943 ] = 8'h00;
    rom[1944 ] = 8'h00;
    rom[1945 ] = 8'h00;
    rom[1946 ] = 8'h00;
    rom[1947 ] = 8'h00;
    rom[1948 ] = 8'h00;
    rom[1949 ] = 8'h00;
    rom[1950 ] = 8'h00;
    rom[1951 ] = 8'h00;
    rom[1952 ] = 8'h00;
    rom[1953 ] = 8'h01;
    rom[1954 ] = 8'h01;
    rom[1955 ] = 8'h01;
    rom[1956 ] = 8'h01;
    rom[1957 ] = 8'h01;
    rom[1958 ] = 8'h07;
    rom[1959 ] = 8'h07;
    rom[1960 ] = 8'h07;
    rom[1961 ] = 8'h1F;
    rom[1962 ] = 8'h1F;
    rom[1963 ] = 8'h1F;
    rom[1964 ] = 8'h1F;
    rom[1965 ] = 8'h1F;
    rom[1966 ] = 8'h1F;
    rom[1967 ] = 8'h1F;
    rom[1968 ] = 8'h1F;
    rom[1969 ] = 8'h1F;
    rom[1970 ] = 8'h1F;
    rom[1971 ] = 8'h1F;
    rom[1972 ] = 8'h1F;
    rom[1973 ] = 8'h1F;
    rom[1974 ] = 8'h1F;
    rom[1975 ] = 8'h1F;
    rom[1976 ] = 8'h1F;
    rom[1977 ] = 8'h1F;
    rom[1978 ] = 8'h1F;
    rom[1979 ] = 8'h1F;
    rom[1980 ] = 8'h1F;
    rom[1981 ] = 8'h1F;
    rom[1982 ] = 8'h1F;
    rom[1983 ] = 8'h1F;
    rom[1984 ] = 8'h1F;
    rom[1985 ] = 8'h1F;
    rom[1986 ] = 8'h1F;
    rom[1987 ] = 8'h1F;
    rom[1988 ] = 8'h1F;
    rom[1989 ] = 8'h1F;
    rom[1990 ] = 8'h07;
    rom[1991 ] = 8'h01;
    rom[1992 ] = 8'h00;
    rom[1993 ] = 8'h00;
    rom[1994 ] = 8'h00;
    rom[1995 ] = 8'h00;
    rom[1996 ] = 8'h00;
    rom[1997 ] = 8'h00;
    rom[1998 ] = 8'h00;
    rom[1999 ] = 8'h00;
    rom[2000 ] = 8'h00;
    rom[2001 ] = 8'h00;
    rom[2002 ] = 8'h00;
    rom[2003 ] = 8'h00;
    rom[2004 ] = 8'h00;
    rom[2005 ] = 8'h00;
    rom[2006 ] = 8'h00;
    rom[2007 ] = 8'h00;
    rom[2008 ] = 8'h00;
    rom[2009 ] = 8'h00;
    rom[2010 ] = 8'h00;
    rom[2011 ] = 8'h00;
    rom[2012 ] = 8'h00;
    rom[2013 ] = 8'h00;
    rom[2014 ] = 8'h00;
    rom[2015 ] = 8'h00;
    rom[2016 ] = 8'h00;
    rom[2017 ] = 8'h00;
    rom[2018 ] = 8'h00;
    rom[2019 ] = 8'h00;
    rom[2020 ] = 8'h00;
    rom[2021 ] = 8'h00;
    rom[2022 ] = 8'h00;
    rom[2023 ] = 8'h00;
    rom[2024 ] = 8'h00;
    rom[2025 ] = 8'h00;
    rom[2026 ] = 8'h00;
    rom[2027 ] = 8'h00;
    rom[2028 ] = 8'h00;
    rom[2029 ] = 8'h00;
    rom[2030 ] = 8'h00;
    rom[2031 ] = 8'h00;
    rom[2032 ] = 8'h00;
    rom[2033 ] = 8'h00;
    rom[2034 ] = 8'h00;
    rom[2035 ] = 8'h00;
    rom[2036 ] = 8'h00;
    rom[2037 ] = 8'h00;
    rom[2038 ] = 8'h00;
    rom[2039 ] = 8'h00;
    rom[2040 ] = 8'h00;
    rom[2041 ] = 8'h00;
    rom[2042 ] = 8'h00;
    rom[2043 ] = 8'h00;
    rom[2044 ] = 8'h00;
    rom[2045 ] = 8'h00;
    rom[2046 ] = 8'h00;
    rom[2047 ] = 8'h00;
end
endmodule
